netcdf elev1 {
dimensions:
	lat = 15 ;
	lon = 10 ;
variables:
	float lat(lat) ;
		lat:name = "latitude" ;
	float lon(lon) ;
		lon:name = "longitude" ;
	short elev(lat, lon) ;
		elev:name = "height" ;
data:
    lat = 6.5, 5.5, 4.5, 3.5, 4.5, 2.5, 1.5, 0.5, -0.5, -1.5, -2.5, -3.5, -4.5, -5.5, -6.5 ;
    lon = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5 ;
}