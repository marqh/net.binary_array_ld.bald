netcdf identity {
    dimensions:
        d0 = 1 ;
        d1 = 1 ;
    variables:
        int var0 ;
        int var1 ;
        int prefix_list ;
            prefix_list:bald__ = "https://www.opengis.net/def/binary-array-ld/";
            prefix_list:skos__ = "http://www.w3.org/2004/02/skos/core#";

    :bald__isPrefixedBy = "prefix_list";
}